`timescale 1 ns/100 ps
// Version: 2022.2 2022.2.0.10


module PF_INIT_MONITOR_C0_PF_INIT_MONITOR_C0_0_PF_INIT_MONITOR(
       FABRIC_POR_N,
       PCIE_INIT_DONE,
       SRAM_INIT_DONE,
       DEVICE_INIT_DONE,
       USRAM_INIT_DONE,
       XCVR_INIT_DONE,
       USRAM_INIT_FROM_SNVM_DONE,
       USRAM_INIT_FROM_UPROM_DONE,
       USRAM_INIT_FROM_SPI_DONE,
       SRAM_INIT_FROM_SNVM_DONE,
       SRAM_INIT_FROM_UPROM_DONE,
       SRAM_INIT_FROM_SPI_DONE,
       AUTOCALIB_DONE,
       BANK_0_VDDI_STATUS,
       BANK_1_VDDI_STATUS,
       BANK_2_VDDI_STATUS,
       BANK_4_VDDI_STATUS,
       BANK_5_VDDI_STATUS,
       BANK_6_VDDI_STATUS,
       BANK_7_VDDI_STATUS
    );
output FABRIC_POR_N;
output PCIE_INIT_DONE;
output SRAM_INIT_DONE;
output DEVICE_INIT_DONE;
output USRAM_INIT_DONE;
output XCVR_INIT_DONE;
output USRAM_INIT_FROM_SNVM_DONE;
output USRAM_INIT_FROM_UPROM_DONE;
output USRAM_INIT_FROM_SPI_DONE;
output SRAM_INIT_FROM_SNVM_DONE;
output SRAM_INIT_FROM_UPROM_DONE;
output SRAM_INIT_FROM_SPI_DONE;
output AUTOCALIB_DONE;
output BANK_0_VDDI_STATUS;
output BANK_1_VDDI_STATUS;
output BANK_2_VDDI_STATUS;
output BANK_4_VDDI_STATUS;
output BANK_5_VDDI_STATUS;
output BANK_6_VDDI_STATUS;
output BANK_7_VDDI_STATUS;

    wire GND_net, VCC_net;
    
    INIT #( .FABRIC_POR_N_SIMULATION_DELAY(1000), .PCIE_INIT_DONE_SIMULATION_DELAY(4000)
        , .SRAM_INIT_DONE_SIMULATION_DELAY(6000), .UIC_INIT_DONE_SIMULATION_DELAY(7000)
        , .USRAM_INIT_DONE_SIMULATION_DELAY(5000) )  I_INIT (
        .FABRIC_POR_N(FABRIC_POR_N), .GPIO_ACTIVE(), .HSIO_ACTIVE(), 
        .PCIE_INIT_DONE(PCIE_INIT_DONE), .RFU({AUTOCALIB_DONE, nc0, 
        nc1, nc2, nc3, SRAM_INIT_FROM_SPI_DONE, 
        SRAM_INIT_FROM_UPROM_DONE, SRAM_INIT_FROM_SNVM_DONE, 
        USRAM_INIT_FROM_SPI_DONE, USRAM_INIT_FROM_UPROM_DONE, 
        USRAM_INIT_FROM_SNVM_DONE, XCVR_INIT_DONE}), .SRAM_INIT_DONE(
        SRAM_INIT_DONE), .UIC_INIT_DONE(DEVICE_INIT_DONE), 
        .USRAM_INIT_DONE(USRAM_INIT_DONE));
    BANKEN #( .BANK_EN_SIMULATION_DELAY(1000), .BANK_NUMBER("bank7")
         )  I_BEN_7 (.BANK_EN(BANK_7_VDDI_STATUS));
    BANKEN #( .BANK_EN_SIMULATION_DELAY(1000), .BANK_NUMBER("bank2")
         )  I_BEN_2 (.BANK_EN(BANK_2_VDDI_STATUS));
    BANKEN #( .BANK_EN_SIMULATION_DELAY(1000), .BANK_NUMBER("bank0")
         )  I_BEN_0 (.BANK_EN(BANK_0_VDDI_STATUS));
    BANKEN #( .BANK_EN_SIMULATION_DELAY(1000), .BANK_NUMBER("bank6")
         )  I_BEN_6 (.BANK_EN(BANK_6_VDDI_STATUS));
    BANKEN #( .BANK_EN_SIMULATION_DELAY(1000), .BANK_NUMBER("bank1")
         )  I_BEN_1 (.BANK_EN(BANK_1_VDDI_STATUS));
    VCC vcc_inst (.Y(VCC_net));
    BANKEN #( .BANK_EN_SIMULATION_DELAY(1000), .BANK_NUMBER("bank5")
         )  I_BEN_5 (.BANK_EN(BANK_5_VDDI_STATUS));
    GND gnd_inst (.Y(GND_net));
    BANKEN #( .BANK_EN_SIMULATION_DELAY(1000), .BANK_NUMBER("bank4")
         )  I_BEN_4 (.BANK_EN(BANK_4_VDDI_STATUS));
    
endmodule
