LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_arith.all;
USE ieee.std_logic_unsigned.all;

package LuSEE_Pkg is


   type Array_7_TO_0   is array (natural range <>)  of STD_LOGIC_VECTOR(7 downto 0);
   type Array_10_TO_0  is array (natural range <>) of STD_LOGIC_VECTOR(10 downto 0);
   type Array_11_TO_0  is array (natural range <>) of STD_LOGIC_VECTOR(11 downto 0);
   type Array_12_TO_0  is array (natural range <>) of STD_LOGIC_VECTOR(12 downto 0);
   type Array_13_TO_0  is array (natural range <>) of STD_LOGIC_VECTOR(13 downto 0);
   type Array_14_TO_0  is array (natural range <>) of STD_LOGIC_VECTOR(14 downto 0);   
   type Array_15_TO_0  is array (natural range <>) of STD_LOGIC_VECTOR(15 downto 0);
   type Array_23_TO_0  is array (natural range <>) of STD_LOGIC_VECTOR(23 downto 0);
   type Array_29_TO_0  is array (natural range <>) of STD_LOGIC_VECTOR(29 downto 0);
     
   
end package;

package body LuSEE_Pkg is

   

end package body LuSEE_Pkg;